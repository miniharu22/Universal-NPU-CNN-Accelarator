`timescale 1ns/10ps

module tb_PE;

	reg clk, reset;

    reg [8*9-1:0] mat_in [0:63];
	reg [8-1:0] weight[0:8];
    reg [8-1:0] mat_out [0:63];

    reg [8-1:0] p_out;
	
	reg [8*9-1:0] in;
	wire [8*9-1:0] weightin;
	wire [8-1:0] out;
	reg en;
	wire out_en;
	
	assign weightin = {weight[0], weight[1], weight[2], weight[3], weight[4], weight[5], weight[6], weight[7], weight[8]}; 

	PE_m P0(in, weightin, 16'b0000_0000_0000_0000, 3'b000, 3'b000, en, out, out_en, clk, reset);
	
	initial
	begin
		clk = 1;
		reset = 0;
		en = 0;
		#12
		reset = 1;
	end
	
	always #5 clk = ~clk;
	
    integer i=0, j=0;

	initial
	begin		
		$readmemh("C://MY/Vivado/UniNPU/UniNPU.srcs/data/input_pe.txt", mat_in);
		$readmemh("C://MY/Vivado/UniNPU/UniNPU.srcs/data/input_pe_wi.txt", weight);
		begin
			#(21);
			for (i=0; i<64; i=i+1)
			begin
				in = mat_in[i];
				en = 1;
				#(10);
			end
		end
	end

	
	integer err = 0;
	initial
	begin		
		$readmemh("C://MY/Vivado/UniNPU/UniNPU.srcs/data/output_pe.txt", mat_out);
		begin
			#(40);    
			for (j=0; j<64; j=j+1)
			begin
                p_out = mat_out[j];
                #(9);
				if (out != p_out) err = err + 1;
				#(1);
			end
		end
	end

endmodule
